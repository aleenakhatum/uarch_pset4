module writeback_stage(
    input wire [6:0] ctrl_in,
    output wire [6:0] ctrl_out
);
    assign ctrl_out = ctrl_in;

endmodule